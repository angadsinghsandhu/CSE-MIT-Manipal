/******************************************************************************

                        #1 : Hello World in Verolog

*******************************************************************************/

module hello_world ;

initial begin
  $display ("Hello World by Angad");
   #10  $finish;
end

endmodule // End of Module hello_world